module circuito_simples (A, B, Y);
input A, B;
output Y;
and AND1 (Y, A, B);
endmodule